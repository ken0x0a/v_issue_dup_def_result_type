module def

pub struct Result<T> {
	data T
	a    string
	b    int
}

pub struct Inner {
	a string
	b int
}

pub struct Inner2 {
	a string
	b int
}

pub struct Inner3 {
	a string
	b int
}
